--	PROCESS (letter)
--	BEGIN
--	CASE letter IS
--		WHEN 'A' => display_code <= "1101001";
--		WHEN 'L' => display_code <= "1101001";
--		WHEN 'T' => display_code <= "1101001";
--		WHEN 'U' => display_code <= "1101001";
--		WHEN 'R' => display_code <= "1101001";
--		WHEN 'C' => display_code <= "1101001";
--		WHEN 'O' => display_code <= "1101001";
--		WHEN '-' => display_code <= "0000000"; 
--	END CASE;

--	CASE num IS
--		WHEN 0 => display_code:= "1000000"; -- nr 0
--		WHEN 1 => display_code:= "1111001"; -- nr 1
--		WHEN 2 => display_code:= "0100100"; -- nr 2
--		WHEN 3 => display_code:= "0110000"; -- nr 3
--		WHEN 4 => display_code:= "0011001"; -- nr 4
--		WHEN 5 => display_code:= "0010010"; -- nr 5
--		WHEN 6 => display_code:= "0000010"; -- nr 6
--		WHEN 7 => display_code:= "1111000"; -- nr 7
--		WHEN 8 => display_code:= "0000000"; -- nr 8
--		WHEN 9 => display_code:= "0011000"; -- nr 9
--		WHEN 0 => display_code:= "1111111"; -- tudo apagado				
--	END CASE;
			



--	END PROCESS;


		