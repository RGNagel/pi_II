--	PROCESS (letter)
--	BEGIN
--	CASE letter IS
--		WHEN 'A' => display_code <= "1101001";
--		WHEN 'L' => display_code <= "1101001";
--		WHEN 'T' => display_code <= "1101001";
--		WHEN 'U' => display_code <= "1101001";
--		WHEN 'R' => display_code <= "1101001";
--		WHEN 'C' => display_code <= "1101001";
--		WHEN 'O' => display_code <= "1101001";
--		WHEN '-' => display_code <= "0000000"; 
--	END CASE;
--	END PROCESS;