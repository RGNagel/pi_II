-- ENTITY FOR CLICK SENSIBILITY

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity setDisplaysNum is
	Port (
		  NUM: IN std_logic_vector ()
   );
end setDisplaysNum;